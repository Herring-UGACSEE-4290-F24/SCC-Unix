module ID();

    

endmodule