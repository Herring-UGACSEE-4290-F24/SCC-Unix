module ID();

    input [31:0] instruction;

    
    

endmodule