module ID();

    input instruction;

    reg [1:0] 1LD;
    reg S;
    reg [3:0] 2LD;
    reg [2:0] ALU_OC; 
    

endmodule