`timescale 1ns/1ns

module DM_tb()

endmodule